module DOL(
  input [63:0] AWDATA);
endmodule
